LIBRARY ieee
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

ENTITY KEYBOARD IS
PORT(
	lin IN : 
)