LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY trans2 IS
PORT(
	clk : IN std_logic;
	rfk : IN std_logic_vector(3 DOWNTO 0);--read from keyboard
	wtk : IN std_logic_vector(3 DOWNTO 0);--read from trans 
	outpu : OUT std_logic_vector (3 DOWNTO 0)
);
END trans2;

ARCHITECTURE behave OF trans2 IS
	SIGNAL buff : std_logic_vector(3 DOWNTO 0);
BEGIN
	outpu <= buff;
	PROCESS(clk)
	BEGIN
		IF(clk'EVENT AND clk = '1') THEN
			CASE rfk & wtk IS
				WHEN "11101110" => buff <= "0001";--1
				WHEN "11101101" => buff <= "0010";--2
				WHEN "11101011" => buff <= "0011";--3
				WHEN "11100111" => buff <= "1010";--a
				WHEN "11011110" => buff <= "0100";--4
				WHEN "11011101" => buff <= "0101";--5
				WHEN "11011011" => buff <= "0110";--6
				WHEN "11010111" => buff <= "1011";--b
				WHEN "10111110" => buff <= "0111";--7
				WHEN "10111101" => buff <= "1000";--8
				WHEN "10111011" => buff <= "1001";--9
				WHEN "10110111" => buff <= "1100";--c
				WHEN "01111110" => buff <= "1110";--e
				WHEN "01111101" => buff <= "0000";--0
				WHEN "01111011" => buff <= "1111";--f
				WHEN "01110111" => buff <= "1101";--d
				WHEN others => null;
			END CASE;
		END IF;
	END PROCESS;
END behave;